pll_10mhz_inst : pll_10mhz PORT MAP (
		inclk0	 => inclk0_sig,
		c0	 => c0_sig
	);
